module Mem (
	input clk,
	input rst,
	input 
);
	
endmodule